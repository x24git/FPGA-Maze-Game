`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    11:09:38 03/09/2018 
// Design Name: 
// Module Name:    maze_selector 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module maze_selector(
    input [7:0] sel,
    input send,
    output reg [maze_flat:0] maze,
    output reg [maze_player_dim:0] player_start,
    output reg [maze_player_dim:0] player_end
    );
`include "maze_parameters.v"	 
reg [maze_player_dim_split:0] index_i;
reg [maze_player_dim_split:0] index_j; 

	 
reg [maze_flat:0] maze_flat_1 = 0;	 
wire [19:0] maze_1[19:0]= {
	20'b10111111111111111111,
	20'b10000001000000101011,
	20'b11111101111110101011,
	20'b10000101000010000001,
	20'b11110001011010101101,
	20'b10010101001010101001,
	20'b11011101011111101011,
	20'b10000001000011000101,
	20'b10111111111100011101,
	20'b10000000000001011101,
	20'b11111101111111000001,
	20'b10000000010000011101,
	20'b11011101000111111001,
	20'b10100001010100000011,
	20'b10001101110001111111,
	20'b11110001000101000001,
	20'b10000100011000010111,
	20'b11110111000010100001,
	20'b10000001000010001101,
	20'b11111111111111111101};
reg[maze_player_dim:0] player_start_1 = 10'b0000100000;
reg[maze_player_dim:0] player_end_1 = 10'b1001010011;

reg [maze_flat:0] maze_flat_2 = 0;	 
wire [19:0] maze_2[19:0]= {
20'b11111111111111111111,
20'b00001000000000000011,
20'b11101110111111111101,
20'b10001010001000001001,
20'b10111010101011111101,
20'b10100010101000001001,
20'b10101111101011111011,
20'b10001000100010001001,
20'b10111110101110111111,
20'b10100000001000001001,
20'b10101011101011101101,
20'b10001010001010100001,
20'b11111111101110101111,
20'b10000000001000000001,
20'b10111110101110111011,
20'b10101000100000001001,
20'b11101011111011101011,
20'b10001000001000101001,
20'b10101111101011100000,
20'b11111111111111111111};

reg[maze_player_dim:0] player_start_2 = 10'b0000000001;
reg[maze_player_dim:0] player_end_2 = 10'b1001110010;

reg [maze_flat:0] maze_flat_3 = 0;	 
wire [19:0] maze_3[19:0]= {
20'b11111111111111111111,
20'b00000000000000100011,
20'b11101110111111111011,
20'b10001000000000100011,
20'b11111011111010101111,
20'b10000010101010001011,
20'b10101110101110111011,
20'b10100010000010001001,
20'b11111010101111101011,
20'b10000000100010000011,
20'b10101110101111111111,
20'b10100010100000000011,
20'b11101110111110111011,
20'b10100010001000001001,
20'b10101011101111101111,
20'b10001010100000100001,
20'b10111010101110101011,
20'b10101000100010101011,
20'b10101011111010101000,
20'b11111111111111111111};

reg[maze_player_dim:0] player_start_3 = 10'b0000000001;
reg[maze_player_dim:0] player_end_3 = 10'b1001110010;

reg [maze_flat:0] maze_flat_4 = 0;	 
wire [19:0] maze_4[19:0]= {
20'b11111111111111111111,
20'b00000000100010001001,
20'b10111110101011101101,
20'b10001010101000001001,
20'b10111010111011101011,
20'b10100000101010000011,
20'b10111011101011101111,
20'b10100000100010101001,
20'b10101011101110111011,
20'b10101010100010100011,
20'b11101010111010111011,
20'b10101000100000001011,
20'b10101110111011111011,
20'b10001010001000100001,
20'b11111010111110111011,
20'b10100010000010000011,
20'b10111011111011111011,
20'b10100000000010000111,
20'b10111110111000110000,
20'b11111111111111111111};

reg[maze_player_dim:0] player_start_4 = 10'b0000000001;
reg[maze_player_dim:0] player_end_4 = 10'b1001110010;

reg [maze_flat:0] maze_flat_5 = 0;	 
wire [19:0] maze_5[19:0]= {
20'b11111111111111111111,
20'b00000000100000000001,
20'b11101011101111111011,
20'b10001000100000001011,
20'b10111010111011111011,
20'b10001010100000001001,
20'b11101111101111101011,
20'b10000000001000101011,
20'b10111010111010111011,
20'b10100010001010100011,
20'b10111011111011101111,
20'b10001000100010001111,
20'b10111110101111111111,
20'b10000010001010001011,
20'b10111010111010101011,
20'b10100010000010100011,
20'b11101010111010110111,
20'b10001010001000100011,
20'b11111011101111101000,
20'b11111111111111111111};

reg[maze_player_dim:0] player_start_5 = 10'b0000000001;
reg[maze_player_dim:0] player_end_5 = 10'b1001110010;

reg [maze_flat:0] maze_flat_6 = 0;	 
wire [19:0] maze_6[19:0]= {
20'b11111111111111111111,
20'b00100000000000100001,
20'b10101111101011101111,
20'b10001000101010000011,
20'b11111110101010101011,
20'b10000010001010101001,
20'b10111111111010101011,
20'b10001010100000101001,
20'b10111010101110111111,
20'b10001010001010100001,
20'b11101011111010101101,
20'b10001000100010001001,
20'b10101011101111101011,
20'b10100000101010001011,
20'b11101110101010111111,
20'b10001000101000001001,
20'b11111010101111100011,
20'b10000010001000001001,
20'b11111111101111101100,
20'b11111111111111111111};

reg[maze_player_dim:0] player_start_6 = 10'b0000000001;
reg[maze_player_dim:0] player_end_6 = 10'b1001110010;

reg [maze_flat:0] maze_flat_7 = 0;	 
wire [19:0] maze_7[19:0]= {
20'b11111111111111111111,
20'b00001000000010001001,
20'b10111111101010101011,
20'b10000000001000100011,
20'b11101111101111111011,
20'b10001000101000001011,
20'b10111110101111101011,
20'b10100000100010101001,
20'b11101111111010101111,
20'b10100000000000100011,
20'b10111111101010101111,
20'b10000000101010001011,
20'b11111110111010111011,
20'b10000000100010000011,
20'b10111011101110111111,
20'b10101000001000000001,
20'b10101011111011111111,
20'b10001010000000000011,
20'b11101110111011111000,
20'b11111111111111111111};

reg[maze_player_dim:0] player_start_7 = 10'b0000000001;
reg[maze_player_dim:0] player_end_7 = 10'b1001110010;

reg [maze_flat:0] maze_flat_8 = 0;	 
wire [19:0] maze_8[19:0]= {
20'b11111111111111111111,
20'b00000010000000001001,
20'b10101110111111101011,
20'b10101000101000101001,
20'b10101010101011101011,
20'b10101010101000101011,
20'b10101011101110111111,
20'b10101000001010000001,
20'b10111111101011111011,
20'b10001010001010101001,
20'b10111010111010101011,
20'b10101000101010100011,
20'b10101011101010111011,
20'b10000010100010100011,
20'b11101110101110111011,
20'b10001000000000001001,
20'b10111011101111101101,
20'b10101010100010000001,
20'b10101010111011111100,
20'b11111111111111111111};

reg[maze_player_dim:0] player_start_8 = 10'b0000000001;
reg[maze_player_dim:0] player_end_8 = 10'b1001110010;

reg [maze_flat:0] maze_flat_default = 0;	 
wire [19:0] maze_default[19:0]= {
	20'b11111111111111111111,
	20'b10000000000000000001,
	20'b10000000000000000001,
	20'b10000000000000000001,
	20'b10000000000000000001,
	20'b10000000000000000001,
	20'b10000000000000000001,
	20'b10000000000000000001,
	20'b10000000000000000001,
	20'b10000000000000000001,
	20'b10000000000000000001,
	20'b10000000000000000001,
	20'b10000000000000000001,
	20'b10000000000000000001,
	20'b10000000000000000001,
	20'b10000000000000000001,
	20'b10000000000000000001,
	20'b10000000000000000001,
	20'b10000000000000000001,	
	20'b11111111111111111111};
reg[maze_player_dim:0] player_start_default = 10'b0100101001;
reg[maze_player_dim:0] player_end_default = 10'b0100101000;
	
	
	
	
always @* begin
	for (index_i = 0; index_i < maze_width; index_i = index_i +1) begin
					for (index_j = 0; index_j < maze_height; index_j = index_j +1) begin
						maze_flat_1[index_i*maze_width+index_j] = maze_1[index_i][index_j];
						maze_flat_2[index_i*maze_width+index_j] = maze_2[index_i][index_j];
						maze_flat_3[index_i*maze_width+index_j] = maze_3[index_i][index_j];
						maze_flat_4[index_i*maze_width+index_j] = maze_4[index_i][index_j];
						maze_flat_5[index_i*maze_width+index_j] = maze_5[index_i][index_j];
						maze_flat_6[index_i*maze_width+index_j] = maze_6[index_i][index_j];
						maze_flat_7[index_i*maze_width+index_j] = maze_7[index_i][index_j];
						maze_flat_8[index_i*maze_width+index_j] = maze_8[index_i][index_j];
						maze_flat_default[index_i*maze_width+index_j] = maze_default[index_i][index_j];
					end
	end


	case(sel)
		8'b00000001: player_start = player_start_1;
		8'b00000010: player_start = player_start_2;
		8'b00000100: player_start = player_start_3;
		8'b00001000: player_start = player_start_4;
		8'b00010000: player_start = player_start_5;
		8'b00100000: player_start = player_start_6;
		8'b01000000: player_start = player_start_7;
		8'b10000000: player_start = player_start_8;
		default: player_start = player_start_default;
	endcase
end

always @(posedge send)begin

	case(sel)
		8'b00000001:begin
			maze = maze_flat_1;
			player_end = player_end_1;
		end
		8'b00000010:begin
			maze = maze_flat_2;
			player_end = player_end_2;
		end
		8'b00000100:begin
			maze = maze_flat_3;
			player_end = player_end_3;
		end
		8'b00001000:begin
			maze = maze_flat_4;
			player_end = player_end_4;
		end
		8'b00010000:begin
			maze = maze_flat_5;
			player_end = player_end_5;
		end
		8'b00100000:begin
			maze = maze_flat_6;
			player_end = player_end_6;
		end
		8'b01000000:begin
			maze = maze_flat_7;
			player_end = player_end_7;
		end
		8'b10000000:begin
			maze = maze_flat_8;
			player_end = player_end_8;
		end
		default: begin
			maze = maze_flat_default;
			player_end = player_end_default;
		end
	endcase
		
end
endmodule
